


module uart
  (
   input        i_Clock,
   input        i_Rx_Serial,
   output       o_Tx_Active,
   output reg   o_Tx_Serial,
   output       o_Tx_Done
   );
	
  parameter c_CLKS_PER_BIT    = 5208;
   
  reg r_Tx_DV = 0;
  wire w_Tx_Done;
  wire w_Tx_Serial;
  wire w_Rx_Done;
  reg [7:0] r_Tx_Byte = 0;
  wire [7:0] w_Rx_Byte;
   
   
  uart_receiver #(.CLKS_PER_BIT(c_CLKS_PER_BIT)) UART_RX_INST
    (.i_Clock(i_Clock),
     .i_Rx_Serial(i_Rx_Serial),
     .o_Rx_DV(w_Rx_Done),
     .o_Rx_Byte(w_Rx_Byte)
     );
   
  uart_transmitter #(.CLKS_PER_BIT(c_CLKS_PER_BIT)) UART_TX_INST
    (.i_Clock(i_Clock),
     .i_Tx_DV(r_Tx_DV),
     .i_Tx_Byte(r_Tx_Byte),
     .o_Tx_Active(o_Tx_Active),
     .o_Tx_Serial(w_Tx_Serial),
     .o_Tx_Done(w_Tx_Done)
     );
 
   
  // Main Testing:
  initial
    begin
       
		o_Tx_Serial <= w_Tx_Serial;
      @(posedge i_Clock);
      @(posedge w_Rx_Done);
      r_Tx_Byte <= w_Rx_Byte;
      @(posedge i_Clock);
      r_Tx_DV <= 1'b1;
		@(posedge i_Clock);
      r_Tx_DV <= 1'b0;
      @(posedge w_Tx_Done);
       
      $display(r_Tx_Byte);
       
    end
   
	assign o_Tx_Done = w_Tx_Done;
endmodule